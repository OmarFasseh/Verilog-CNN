//test bench for floating-point multiplication
module mul_flp_tb;

parameter EXPONENT_WIDTH = 8;
parameter MANTISSA_WIDTH = 23;

reg [31:0] flp_a, flp_b;
reg clock;
wire sign;
wire [7:0] exponent;
wire [8:0] exp_sum;
wire [22:0] prod;
initial
begin
clock = 1;

//+5 x +3 = +15
// s ----e---- --------------f-------------
#2 flp_a = 32'b01000000101000000000000000000000;
flp_b = 32'b01000000010000000000000000000000;
//+6 x +4 = +24
// s ----e---- --------------f-------------
#2 flp_a = 32'b01000000110000000000000000000000;
flp_b = 32'b01000000100000000000000000000000;
//-5 x +5 = -25
// s ----e---- --------------f-------------
#2 flp_a = 32'b11000000101000000000000000000000;
flp_b = 32'b01000000101000000000000000000000;
//+7 x -5 = -35
// s ----e---- --------------f-------------
#2 flp_a = 32'b01000000111000000000000000000000;
flp_b = 32'b11000000101000000000000000000000;
//+25 x +25 = +625
// s ----e---- --------------f-------------
#2 flp_a = 32'b01000001110010000000000000000000;
flp_b = 32'b01000001110010000000000000000000;
//continued on next page

//+76 x +55 = +4180
// s ----e---- --------------f-------------
#2 flp_a = 32'b01000010100110000000000000000000;
flp_b = 32'b01000010010111000000000000000000;
//-48 x -17 = +816
// s ----e---- --------------f-------------
#2 flp_a = 32'b11000010010000000000000000000000;
flp_b = 32'b11000001100010000000000000000000;
//+3724 x +853 = +3,176,572
// s ----e---- --------------f-------------
#2 flp_a = 32'b01000101011010001100000000000000;
flp_b = 32'b01000100010101010100000000000000;

//+5 * 0.00381924584508 = 0.0.01909622922;
#2 flp_a = 32'b01000000101000000000000000000000;
flp_b = 32'b00111011011110100100110001010000;

//More TESTS
#2
flp_a= 32'b00000000000000000000000000000000; //0  
flp_b= 32'b00000000000000000000000000000000; //0  

#2

flp_a= 32'b11000000111100000000000000000000; //-7.5  
flp_b= 32'b01000010000011000000000000000000; //35   

#2

flp_a= 32'b01000010001101000000000000000000; //45  
flp_b= 32'b11000000010000000000000000000000; //-3   

#2

flp_a= 32'b01000000000000000000000000000000; //2  
flp_b= 32'b01000000011000000000000000000000; //3.5   


#2

flp_a= 32'b01000001000100000000000000000000; //9  
flp_b= 32'b11000010101100000000000000000000; //-88  


#2

flp_a= 32'b00000000000000000000000000000000; //0  
flp_b= 32'b01000001010000000000000000000000; //12  

#2

flp_a =32'b00111111000000000000000000000000; //.5  
flp_b =32'b00111111000000000000000000000000; //.5  

#2

flp_a =32'b11000010110001100000000000000000; //-99  
flp_b =32'b11000010000001000000000000000000; //-33  

#2

flp_a =32'b00111111000000000000000000000000; //0.5  
flp_b =32'b00111110100110011001100110011000; //0.3  


#2

flp_a =32'b00111110010011001100110011001100; //0.2  
flp_b =32'b00111111000000000000000000000000; //0.5  

#2

flp_a =32'b01000000001000000000000000000000; //2.5  
flp_b =32'b01000000100100000000000000000000; //4.5  

#2

flp_a =32'b01000000001000000000000000000000; //2.5  
flp_b =32'b01000001001000000000000000000000; //10  
#2 $stop;
end


always begin
     #1  clock = ~clock; 
    end
        
//instantiate the module into the test bench
fpMul #(.EXPONENT_WIDTH(EXPONENT_WIDTH), .MANTISSA_WIDTH(MANTISSA_WIDTH)) inst1 (
.flp_a(flp_a),
.flp_b(flp_b),
.sign(sign),
.exponent(exponent),
.prod(prod),
.clk(clock)
);
endmodule
