//test bench for floating-point addition
`timescale 1ns / 1ps

module add_flp3_tb;

parameter EXPONENT_WIDTH = 5;
parameter MANTISSA_WIDTH = 10;
    reg [EXPONENT_WIDTH+MANTISSA_WIDTH:0] A, B;
    reg clock;
    wire sign_C;
    wire [EXPONENT_WIDTH-1:0] exp_C;
    wire [MANTISSA_WIDTH-1:0] mantissa_C;
    initial //display variables
    $monitor ("sign=%b, exp_biased=%b, sum=%b",sign_C, exp_C, mantissa_C);
    
    initial //apply input vectors
    begin
        clock = 1;
        //+7.25 + + 0.375 = + 7.625 = 0b0100011110100000
                // s ----e---- --------------M-------------
        #2 A = 32'b0100011101000000;
           B = 32'b0011011000000000;
        //+6 + +7 = + 13 = 0b0100101010000000
                // s ----e---- --------------M-------------
        #2 A = 32'b0100011000000000;
           B = 32'b0100011100000000;
        // -7 + -3 = -10 = 0b1100100100000000
        #2 A = 32'b1100011100000000;
           B = 32'b1100001000000000;
        // 7 + -3 = 4 = 0b0100010000000000
        #2 A = 32'b0100011100000000;
           B = 32'b1100001000000000;
        // -7.0 + 3 = -4 = 0b1100010000000000
        #2 A = 32'b1100011100000000;
           B = 32'b0100001000000000; 
        //65 - 63 = 2 = 0b0100000000000000
        #2 A = 32'b0101010000010000;
           B = 32'b1101001111100000;
           //4 - 4 = 0 = 0b0000000000000000
        #2 A = 32'b0100010000000000;
           B = 32'b0100010000000000;
         #2
           //MOAZ TEST CASES for 32 bit, remove later:
        /*A= 32'b00000000000000000000000000000000; //0 dec
        B= 32'b00000000000000000000000000000000; //0 dec

        #2

        A= 32'b11000010000100000000000000000000; //-36 dec
        B= 32'b01000001001000000000000000000000; //10 dec

        #2

        A= 32'b01000001000100000000000000000000; //9 dec
        B= 32'b11000010101100000000000000000000; //-88 dec


        #2

        A= 32'b00000000000000000000000000000000; //0 dec
        B= 32'b01000001010000000000000000000000; //12 dec

        #2

        A =32'b10111111000000000000000000000000; //-0.5dec
        B =32'b00111111000000000000000000000000; //0.5 dec

        #2

        A =32'b11000010110001100000000000000000; //-99 dec
        B =32'b11000010000001000000000000000000; //-33 dec

        #2

        A =32'b00111111000000000000000000000000; //0.5 dec
        B =32'b10111110100110011001100110011000; //-0.3 dec


        #2

        A =32'b00111110010011001100110011001100; //0.2 dec
        B =32'b00111111000000000000000000000000; //0.5 dec

        #2

        A =32'b01000000001000000000000000000000; //2.5 dec
        B =32'b11000000100100000000000000000000; //-4.5 dec

        #2

        A =32'b01000000001000000000000000000000; //2.5 dec
        B =32'b01000001001000000000000000000000; //10 dec       
        #2

        A = 32'b01000000100000000000000000000000; //4
        B = 32'b10111111100000000000000000000000; //-1*/
        #2 $stop;
    end
    
    always begin
         #1  clock = ~clock; 
        end
    
    fp_add_2 #(.EXPONENT_WIDTH(EXPONENT_WIDTH), .MANTISSA_WIDTH(MANTISSA_WIDTH))
    fp_add1 ( //instantiate the module
    .A_FP(A),
    .B_FP(B),
    .sign(sign_C),
    .exponent(exp_C),
    .mantissa(mantissa_C),
    .clk(clock));
endmodule
